Adm Circuit

;in1 and in2 are input ports, out1 and out2 are output ports

M1 N015 in1 N018 N018 CMOSN l=0.8u w=399.0422985u
M3 N009 N013 N011 N011 CMOSN l=0.8u w=3.832402235u
M4 N009 N008 N006 N006 CMOSP l=0.8u w=0.08726248081u
M5 N006 N005 N003 N003 CMOSP l=0.8u w=0.08726248081u
M8 N005 N005 N002 N002 CMOSP l=0.8u w=87.26248481u
M9 N008 N008 N005 N005 CMOSP l=0.8u w=87.26248481u
M10 N013 N013 N014 N014 CMOSN l=0.8u w=3832.402235u
I1 N008 N013 50�
V1 in1 in2 SINE(0 10m 1k) AC 10m
V2 in2 0 124.7m
V3 N001 0 3.5
M2 N011 N014 N015 N015 CMOSN l=0.8u w=3.832402235u
M11 N014 N014 N017 N017 CMOSN l=0.8u w=977.5538809u
M7 N002 N002 N001 N001 CMOSP l=0.8u w=319.4316672u
M6 N003 N002 N001 N001 CMOSP l=0.8u w=0.3194316472u
M12 N016 in2 N018 N018 CMOSN l=0.8u w=399.0422985u
M14 N010 N013 N012 N012 CMOSN l=0.8u w=3.832402235u
M15 N010 N008 N007 N007 CMOSP l=0.8u w=0.08726248481u
M16 N007 N005 N004 N004 CMOSP l=0.8u w=0.08726248481u
M13 N012 N014 N016 N016 CMOSN l=0.8u w=3.832402235u
M17 N004 N002 N001 N001 CMOSP l=0.8u w=0.3194316472u
M18 N018 N017 N020 N020 CMOSN l=0.8u w=3.547042653u
M19 N020 N019 0 0 CMOSN l=0.8u w=3.547042653u
M20 N017 N017 N019 N019 CMOSN l=0.8u w=1773.521327u
M21 N019 N019 0 0 CMOSN l=0.8u w=1773.521327u
C1 out1 N009 1p
C2 N010 out2 1p

.ac dec 100 1 1G

.lib mosis_350.lib

.end
